��72      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby_wsp��wzrost��leki�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh&hNhJ�
hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h4�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh(�scalar���hJC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hK�
node_count�K	�nodes�h*h-K ��h/��R�(KK	��h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h{h4�i8�����R�(KhKNNNJ����J����K t�bK ��h|h�K��h}h�K��h~h[K��hh[K ��h�h�K(��h�h[K0��uK8KKt�b�B�                             N@�q�q��?             H@                           @p9W��S�?             C@                          �E@     ��?             @@������������������������       �z�G�z�?             4@������������������������       ��q�q�?             (@������������������������       �                     @                          @h@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�t�b�values�h*h-K ��h/��R�(KK	KK��h[�C�      3@      =@      &@      ;@      &@      5@      @      0@      @      @              @       @       @       @                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ/��hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                             h@�q�q�?!             H@                          �E@�q�q�?            �C@                          Pd@8�Z$���?
             *@������������������������       �                     �?������������������������       ��8��8��?	             (@                            @$�q-�?             :@������������������������       �                     7@������������������������       ��q�q�?             @	                           �?�<ݚ�?             "@
                         yJ@@�q�q�?             @������������������������       �                     �?������������������������       �      �?              @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      <@      4@      :@      *@       @      &@      �?              �?      &@      8@       @      7@              �?       @       @      @       @      �?      �?              �?      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJu�7hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            @K@�q���?             H@                           @�c�Α�?             =@                         ��g@���Q��?             $@������������������������       �                     @������������������������       �z�G�z�?             @                          �E@�KM�]�?             3@������������������������       �      �?	             0@������������������������       ��q�q�?             @	       
                  �%g@�KM�]�?	             3@������������������������       �                     (@                            @����X�?             @������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      9@      7@       @      5@      @      @      @              �?      @       @      1@      �?      .@      �?       @      1@       @      (@              @       @      @                       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��!XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrK	hsh*h-K ��h/��R�(KK	��hz�B�                              �?�q���?             H@������������������������       �                     &@                         �%g@؀�:M�?            �B@                           �?����X�?             ,@������������������������       �z�G�z�?             @������������������������       �                     "@                          �h@�㙢�c�?             7@������������������������       ����y4F�?             3@������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK	KK��h[�C�      9@      7@      &@              ,@      7@      $@      @      �?      @      "@              @      3@      @      .@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJC�NhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                             @      �?#             H@                         �%g@�5��?             ;@                          �:@@4և���?
             ,@������������������������       ��q�q�?             @������������������������       �                     &@                            @�θ�?
             *@������������������������       �      �?              @������������������������       �                     @	                          �M@�ՙ/�?             5@
                            @�E��ӭ�?             2@������������������������       ��eP*L��?	             &@������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      8@      8@      0@      &@      *@      �?       @      �?      &@              @      $@      @      @              @       @      *@      @      *@      @      @              @      @        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�R�[hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            �E@      �?             H@                          Pd@�+e�X�?             9@������������������������       �                      @                          �<@�㙢�c�?             7@������������������������       �                     "@������������������������       �����X�?             ,@       
                     @��<b���?             7@       	                   �g@�KM�]�?             3@������������������������       �        
             1@������������������������       �                      @                           R@      �?             @������������������������       �                     �?������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      8@      8@      @      3@       @              @      3@              "@      @      $@      2@      @      1@       @      1@                       @      �?      @      �?                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�v}hG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                            �E@r�qG�?             H@                           0@p�ݯ��?             3@������������������������       �                     @                         ��e@      �?
             0@������������������������       �                     @������������������������       ��	j*D�?             *@                           �?д>��C�?             =@������������������������       �                     .@	       
                  y
F@X�Cc�?
             ,@������������������������       �                     @������������������������       �X�<ݚ�?             "@�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      ?@      1@      @      (@      @              @      (@              @      @      "@      8@      @      .@              "@      @      @              @      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJg}�XhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                            pg@      �?             H@                            @V�a�� �?             =@                            �?      �?             8@������������������������       �                     &@������������������������       ��θ�?             *@                          �d@���Q��?             @������������������������       �                      @������������������������       ��q�q�?             @	       
                  y�H@�}�+r��?             3@������������������������       �                     .@                          `P@      �?             @������������������������       �      �?              @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      8@      8@      7@      @      5@      @      &@              $@      @       @      @               @       @      �?      �?      2@              .@      �?      @      �?      �?               @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ	�tlhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�Bh                              �?      �?             H@                          �g@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @                            @<=�,S��?            �A@                          �E@��
ц��?             :@������������������������       �������?             1@������������������������       ������H�?             "@	       
                   0f@�����H�?             "@������������������������       �      �?              @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      8@      8@      &@       @      &@                       @      *@      6@      (@      ,@      @      *@       @      �?      �?       @      �?      �?              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�ޡhG        hNhG        hAKhBKhCh*h-K ��h/��R�(KK��h[�C              �?�t�bhOh`hJC       ���R�hdKhehhKh*h-K ��h/��R�(KK��hJ�C       �t�bK��R�}�(hKhrKhsh*h-K ��h/��R�(KK��hz�B�                           y�H@r�qG�?             H@                            @r�q��?             8@                          �h@�G��l��?             5@������������������������       �ҳ�wY;�?
             1@������������������������       �                     @������������������������       �                     @       
                    @r�q��?             8@       	                    @�X�<ݺ?             2@������������������������       �ףp=
�?             $@������������������������       �                      @                            @      �?             @������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KKKK��h[�C�      ?@      1@      &@      *@      &@      $@      &@      @              @              @      4@      @      1@      �?      "@      �?       @              @      @      @                      @�t�bubhhubehhub.